// soc_system.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module soc_system (
		output wire         axi_avl_clk_clk,               //       axi_avl_clk.clk
		input  wire         clk_clk,                       //               clk.clk
		input  wire         f2h_sdram0_clock_clk,          //  f2h_sdram0_clock.clk
		input  wire [27:0]  f2h_sdram0_data_address,       //   f2h_sdram0_data.address
		input  wire [7:0]   f2h_sdram0_data_burstcount,    //                  .burstcount
		output wire         f2h_sdram0_data_waitrequest,   //                  .waitrequest
		output wire [127:0] f2h_sdram0_data_readdata,      //                  .readdata
		output wire         f2h_sdram0_data_readdatavalid, //                  .readdatavalid
		input  wire         f2h_sdram0_data_read,          //                  .read
		input  wire [127:0] f2h_sdram0_data_writedata,     //                  .writedata
		input  wire [15:0]  f2h_sdram0_data_byteenable,    //                  .byteenable
		input  wire         f2h_sdram0_data_write,         //                  .write
		output wire         hps_0_h2f_reset_reset_n,       //   hps_0_h2f_reset.reset_n
		input  wire         hps_f2h_axi_clock_clk,         // hps_f2h_axi_clock.clk
		input  wire [7:0]   hps_f2h_axi_slave_awid,        // hps_f2h_axi_slave.awid
		input  wire [31:0]  hps_f2h_axi_slave_awaddr,      //                  .awaddr
		input  wire [3:0]   hps_f2h_axi_slave_awlen,       //                  .awlen
		input  wire [2:0]   hps_f2h_axi_slave_awsize,      //                  .awsize
		input  wire [1:0]   hps_f2h_axi_slave_awburst,     //                  .awburst
		input  wire [1:0]   hps_f2h_axi_slave_awlock,      //                  .awlock
		input  wire [3:0]   hps_f2h_axi_slave_awcache,     //                  .awcache
		input  wire [2:0]   hps_f2h_axi_slave_awprot,      //                  .awprot
		input  wire         hps_f2h_axi_slave_awvalid,     //                  .awvalid
		output wire         hps_f2h_axi_slave_awready,     //                  .awready
		input  wire [4:0]   hps_f2h_axi_slave_awuser,      //                  .awuser
		input  wire [7:0]   hps_f2h_axi_slave_wid,         //                  .wid
		input  wire [31:0]  hps_f2h_axi_slave_wdata,       //                  .wdata
		input  wire [3:0]   hps_f2h_axi_slave_wstrb,       //                  .wstrb
		input  wire         hps_f2h_axi_slave_wlast,       //                  .wlast
		input  wire         hps_f2h_axi_slave_wvalid,      //                  .wvalid
		output wire         hps_f2h_axi_slave_wready,      //                  .wready
		output wire [7:0]   hps_f2h_axi_slave_bid,         //                  .bid
		output wire [1:0]   hps_f2h_axi_slave_bresp,       //                  .bresp
		output wire         hps_f2h_axi_slave_bvalid,      //                  .bvalid
		input  wire         hps_f2h_axi_slave_bready,      //                  .bready
		input  wire [7:0]   hps_f2h_axi_slave_arid,        //                  .arid
		input  wire [31:0]  hps_f2h_axi_slave_araddr,      //                  .araddr
		input  wire [3:0]   hps_f2h_axi_slave_arlen,       //                  .arlen
		input  wire [2:0]   hps_f2h_axi_slave_arsize,      //                  .arsize
		input  wire [1:0]   hps_f2h_axi_slave_arburst,     //                  .arburst
		input  wire [1:0]   hps_f2h_axi_slave_arlock,      //                  .arlock
		input  wire [3:0]   hps_f2h_axi_slave_arcache,     //                  .arcache
		input  wire [2:0]   hps_f2h_axi_slave_arprot,      //                  .arprot
		input  wire         hps_f2h_axi_slave_arvalid,     //                  .arvalid
		output wire         hps_f2h_axi_slave_arready,     //                  .arready
		input  wire [4:0]   hps_f2h_axi_slave_aruser,      //                  .aruser
		output wire [7:0]   hps_f2h_axi_slave_rid,         //                  .rid
		output wire [31:0]  hps_f2h_axi_slave_rdata,       //                  .rdata
		output wire [1:0]   hps_f2h_axi_slave_rresp,       //                  .rresp
		output wire         hps_f2h_axi_slave_rlast,       //                  .rlast
		output wire         hps_f2h_axi_slave_rvalid,      //                  .rvalid
		input  wire         hps_f2h_axi_slave_rready,      //                  .rready
		inout  wire         hps_io_hps_io_sdio_inst_CMD,   //            hps_io.hps_io_sdio_inst_CMD
		inout  wire         hps_io_hps_io_sdio_inst_D0,    //                  .hps_io_sdio_inst_D0
		inout  wire         hps_io_hps_io_sdio_inst_D1,    //                  .hps_io_sdio_inst_D1
		output wire         hps_io_hps_io_sdio_inst_CLK,   //                  .hps_io_sdio_inst_CLK
		inout  wire         hps_io_hps_io_sdio_inst_D2,    //                  .hps_io_sdio_inst_D2
		inout  wire         hps_io_hps_io_sdio_inst_D3,    //                  .hps_io_sdio_inst_D3
		input  wire         hps_io_hps_io_uart0_inst_RX,   //                  .hps_io_uart0_inst_RX
		output wire         hps_io_hps_io_uart0_inst_TX,   //                  .hps_io_uart0_inst_TX
		output wire [14:0]  memory_mem_a,                  //            memory.mem_a
		output wire [2:0]   memory_mem_ba,                 //                  .mem_ba
		output wire         memory_mem_ck,                 //                  .mem_ck
		output wire         memory_mem_ck_n,               //                  .mem_ck_n
		output wire         memory_mem_cke,                //                  .mem_cke
		output wire         memory_mem_cs_n,               //                  .mem_cs_n
		output wire         memory_mem_ras_n,              //                  .mem_ras_n
		output wire         memory_mem_cas_n,              //                  .mem_cas_n
		output wire         memory_mem_we_n,               //                  .mem_we_n
		output wire         memory_mem_reset_n,            //                  .mem_reset_n
		inout  wire [31:0]  memory_mem_dq,                 //                  .mem_dq
		inout  wire [3:0]   memory_mem_dqs,                //                  .mem_dqs
		inout  wire [3:0]   memory_mem_dqs_n,              //                  .mem_dqs_n
		output wire         memory_mem_odt,                //                  .mem_odt
		output wire [3:0]   memory_mem_dm,                 //                  .mem_dm
		input  wire         memory_oct_rzqin,              //                  .oct_rzqin
		output wire         pll_0_locked_export,           //      pll_0_locked.export
		input  wire         reset_reset_n                  //             reset.reset_n
	);

	soc_system_hps_0 #(
		.F2S_Width (1),
		.S2F_Width (0)
	) hps_0 (
		.mem_a                    (memory_mem_a),                  //           memory.mem_a
		.mem_ba                   (memory_mem_ba),                 //                 .mem_ba
		.mem_ck                   (memory_mem_ck),                 //                 .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),               //                 .mem_ck_n
		.mem_cke                  (memory_mem_cke),                //                 .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),               //                 .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),              //                 .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),              //                 .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),               //                 .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),            //                 .mem_reset_n
		.mem_dq                   (memory_mem_dq),                 //                 .mem_dq
		.mem_dqs                  (memory_mem_dqs),                //                 .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),              //                 .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                //                 .mem_odt
		.mem_dm                   (memory_mem_dm),                 //                 .mem_dm
		.oct_rzqin                (memory_oct_rzqin),              //                 .oct_rzqin
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),   //           hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),    //                 .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),    //                 .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),   //                 .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),    //                 .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),    //                 .hps_io_sdio_inst_D3
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),   //                 .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),   //                 .hps_io_uart0_inst_TX
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),       //        h2f_reset.reset_n
		.f2h_sdram0_clk           (f2h_sdram0_clock_clk),          // f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (f2h_sdram0_data_address),       //  f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (f2h_sdram0_data_burstcount),    //                 .burstcount
		.f2h_sdram0_WAITREQUEST   (f2h_sdram0_data_waitrequest),   //                 .waitrequest
		.f2h_sdram0_READDATA      (f2h_sdram0_data_readdata),      //                 .readdata
		.f2h_sdram0_READDATAVALID (f2h_sdram0_data_readdatavalid), //                 .readdatavalid
		.f2h_sdram0_READ          (f2h_sdram0_data_read),          //                 .read
		.f2h_sdram0_WRITEDATA     (f2h_sdram0_data_writedata),     //                 .writedata
		.f2h_sdram0_BYTEENABLE    (f2h_sdram0_data_byteenable),    //                 .byteenable
		.f2h_sdram0_WRITE         (f2h_sdram0_data_write),         //                 .write
		.f2h_axi_clk              (hps_f2h_axi_clock_clk),         //    f2h_axi_clock.clk
		.f2h_AWID                 (hps_f2h_axi_slave_awid),        //    f2h_axi_slave.awid
		.f2h_AWADDR               (hps_f2h_axi_slave_awaddr),      //                 .awaddr
		.f2h_AWLEN                (hps_f2h_axi_slave_awlen),       //                 .awlen
		.f2h_AWSIZE               (hps_f2h_axi_slave_awsize),      //                 .awsize
		.f2h_AWBURST              (hps_f2h_axi_slave_awburst),     //                 .awburst
		.f2h_AWLOCK               (hps_f2h_axi_slave_awlock),      //                 .awlock
		.f2h_AWCACHE              (hps_f2h_axi_slave_awcache),     //                 .awcache
		.f2h_AWPROT               (hps_f2h_axi_slave_awprot),      //                 .awprot
		.f2h_AWVALID              (hps_f2h_axi_slave_awvalid),     //                 .awvalid
		.f2h_AWREADY              (hps_f2h_axi_slave_awready),     //                 .awready
		.f2h_AWUSER               (hps_f2h_axi_slave_awuser),      //                 .awuser
		.f2h_WID                  (hps_f2h_axi_slave_wid),         //                 .wid
		.f2h_WDATA                (hps_f2h_axi_slave_wdata),       //                 .wdata
		.f2h_WSTRB                (hps_f2h_axi_slave_wstrb),       //                 .wstrb
		.f2h_WLAST                (hps_f2h_axi_slave_wlast),       //                 .wlast
		.f2h_WVALID               (hps_f2h_axi_slave_wvalid),      //                 .wvalid
		.f2h_WREADY               (hps_f2h_axi_slave_wready),      //                 .wready
		.f2h_BID                  (hps_f2h_axi_slave_bid),         //                 .bid
		.f2h_BRESP                (hps_f2h_axi_slave_bresp),       //                 .bresp
		.f2h_BVALID               (hps_f2h_axi_slave_bvalid),      //                 .bvalid
		.f2h_BREADY               (hps_f2h_axi_slave_bready),      //                 .bready
		.f2h_ARID                 (hps_f2h_axi_slave_arid),        //                 .arid
		.f2h_ARADDR               (hps_f2h_axi_slave_araddr),      //                 .araddr
		.f2h_ARLEN                (hps_f2h_axi_slave_arlen),       //                 .arlen
		.f2h_ARSIZE               (hps_f2h_axi_slave_arsize),      //                 .arsize
		.f2h_ARBURST              (hps_f2h_axi_slave_arburst),     //                 .arburst
		.f2h_ARLOCK               (hps_f2h_axi_slave_arlock),      //                 .arlock
		.f2h_ARCACHE              (hps_f2h_axi_slave_arcache),     //                 .arcache
		.f2h_ARPROT               (hps_f2h_axi_slave_arprot),      //                 .arprot
		.f2h_ARVALID              (hps_f2h_axi_slave_arvalid),     //                 .arvalid
		.f2h_ARREADY              (hps_f2h_axi_slave_arready),     //                 .arready
		.f2h_ARUSER               (hps_f2h_axi_slave_aruser),      //                 .aruser
		.f2h_RID                  (hps_f2h_axi_slave_rid),         //                 .rid
		.f2h_RDATA                (hps_f2h_axi_slave_rdata),       //                 .rdata
		.f2h_RRESP                (hps_f2h_axi_slave_rresp),       //                 .rresp
		.f2h_RLAST                (hps_f2h_axi_slave_rlast),       //                 .rlast
		.f2h_RVALID               (hps_f2h_axi_slave_rvalid),      //                 .rvalid
		.f2h_RREADY               (hps_f2h_axi_slave_rready)       //                 .rready
	);

	soc_system_pll_0 pll_0 (
		.refclk   (clk_clk),             //  refclk.clk
		.rst      (~reset_reset_n),      //   reset.reset
		.outclk_0 (axi_avl_clk_clk),     // outclk0.clk
		.locked   (pll_0_locked_export)  //  locked.export
	);

endmodule
